library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity control_unit is
    port (
        clock: in std_ulogic;
        reset: in std_ulogic;

        start: in std_ulogic;

        -- Memory Driver Interface
        memory_driver_start: out std_ulogic;
        memory_driver_address: out std_ulogic_vector(23 downto 0);

        memory_driver_data: in std_ulogic_vector(7 downto 0);
        memory_driver_done: in std_ulogic;

        -- Audio Driver Interface
        audio_driver_play: out std_ulogic;
        audio_driver_done: in std_ulogic;

        -- Audio Fifo
        audio_fifo_write_enable: out std_ulogic;
        audio_fifo_data_in: out std_ulogic_vector(7 downto 0);
        audio_fifo_full: in std_ulogic;

        -- Video Driver Interface
        video_driver_play: out std_ulogic;
        video_driver_done: in std_ulogic;

        -- Video Fifo
        video_fifo_write_enable: out std_ulogic;
        video_fifo_data_in: out std_ulogic_vector(7 downto 0);
        video_fifo_full: in std_ulogic
    );
end entity;

architecture arch of control_unit is
    type state_t is (
        IDLE, READ_HEADER, PARSE_HEADER,
        WAIT_FOR_DATA, REQUEST_DATA, WAIT_FOR_EMPTY_SLOT,
        DONE
    );
    signal state, state_next: state_t;

    signal header, header_next: std_ulogic_vector(10 * 8 - 1 downto 0);
    alias signature_begin: std_ulogic_vector(7 downto 0) is header(7 downto 0);
    alias audio_length: std_ulogic_vector(memory_driver_address'range) is header(8 + memory_driver_address'length - 1 downto 8);
    alias video_length: std_ulogic_vector(memory_driver_address'range) is header(8 + 32 + memory_driver_address'length - 1 downto 8 + 32);
    alias signature_end: std_ulogic_vector(7 downto 0) is header(7 + 32 + 32 + 8 downto 32 + 32 + 8);

    signal audio_pointer, audio_pointer_next: std_ulogic_vector(memory_driver_address'range);
    signal audio_end_address, audio_end_address_next: std_ulogic_vector(memory_driver_address'range);

    signal video_pointer, video_pointer_next: std_ulogic_vector(memory_driver_address'range);
    signal video_end_address, video_end_address_next: std_ulogic_vector(memory_driver_address'range);

    -- If this signal is '1', read and wait for audio, if it's '0', read and wait for video.
    signal read_audio_n_video, read_audio_n_video_next: std_ulogic;

    signal start_playback, start_playback_next: std_ulogic;

    signal audio_loaded, audio_loaded_next: std_ulogic;
    signal video_loaded, video_loaded_next: std_ulogic;
begin
    seq: process (clock)
    begin
        if rising_edge(clock) then
            if reset = '1' then
                state <= IDLE;

                header <= (others => '0');

                audio_pointer <= (others => '0');
                audio_end_address <= (others => '0');

                video_pointer <= (others => '0');
                video_end_address <= (others => '0');

                read_audio_n_video <= '1';

                start_playback <= '0';

                audio_loaded <= '0';
                video_loaded <= '0';
            else
                state <= state_next;

                header <= header_next;

                audio_pointer <= audio_pointer_next;
                audio_end_address <= audio_end_address_next;

                video_pointer <= video_pointer_next;
                video_end_address <= video_end_address_next;

                read_audio_n_video <= read_audio_n_video_next;

                start_playback <= start_playback_next;

                audio_loaded <= audio_loaded_next;
                video_loaded <= video_loaded_next;
            end if;
        end if;
    end process;

    fsm: process (
        state, start,
        header, memory_driver_done, memory_driver_data,
        audio_fifo_full, audio_pointer, audio_end_address,
        video_fifo_full, video_pointer, video_end_address,
        read_audio_n_video, start_playback,
        audio_driver_done, video_driver_done,
        audio_loaded, video_loaded
    )
        variable u_audio_pointer, u_video_pointer: unsigned(audio_pointer'range);
        variable u_audio_length, u_video_length: unsigned(audio_length'range);
    begin
        u_audio_pointer := unsigned(audio_pointer);
        u_video_pointer := unsigned(video_pointer);

        u_audio_length := unsigned(audio_length);
        u_video_length := unsigned(video_length);

        state_next <= state;

        header_next <= header;

        audio_fifo_data_in <= (others => '0');
        audio_fifo_write_enable <= '0';

        audio_pointer_next <= audio_pointer;
        audio_end_address_next <= audio_end_address;

        video_fifo_data_in <= (others => '0');
        video_fifo_write_enable <= '0';

        video_pointer_next <= video_pointer;
        video_end_address_next <= video_end_address;

        read_audio_n_video_next <= read_audio_n_video;

        memory_driver_start <= '0';
        memory_driver_address <= (others => '0');

        start_playback_next <= start_playback;

        audio_driver_play <= '0';
        video_driver_play <= '0';

        audio_loaded_next <= audio_loaded;
        video_loaded_next <= video_loaded;

        case state is
            when IDLE =>
                if start = '1' then
                    state_next <= READ_HEADER;

                    -- We are reading the header first, not the audio but instead of spending
                    -- more hardware to have designated flipflops to hold the current address
                    -- of the header, we can simply use the audio pointer.
                    -- This also has the neat effect, that it lands on the first audio byte
                    -- if audio was included!
                    memory_driver_start <= '1';
                    memory_driver_address <= std_ulogic_vector(to_unsigned(0, memory_driver_address'length));

                    -- Advance the audio pointer to the next address.
                    audio_pointer_next <= std_ulogic_vector(to_unsigned(1, audio_pointer_next'length));

                    audio_loaded_next <= '0';
                    video_loaded_next <= '0';

                    start_playback_next <= '0';
                end if;

            when READ_HEADER =>
                if memory_driver_done = '1' then
                    -- Insert from the MSB otherwise the endianness will change.
                    header_next(header'length - 1 downto header'length - memory_driver_data'length) <= memory_driver_data;
                    header_next(header'length - memory_driver_data'length - 1 downto 0) <= header(header'length - 1 downto memory_driver_data'length);

                    -- Since we are reading from IDLE -> READ_HEADER the address was incremented already.
                    -- This means that address contains the next address so we have to check for
                    -- header'length / 8 and not -1.
                    if u_audio_pointer = header'length / 8 then
                        state_next <= PARSE_HEADER;
                    else
                        memory_driver_start <= '1';
                        memory_driver_address <= audio_pointer;

                        audio_pointer_next <= std_ulogic_vector(u_audio_pointer + 1);
                    end if;
                end if;

            when PARSE_HEADER =>
                if unsigned(signature_begin) = to_unsigned(character'pos('A'), 8)
                    and unsigned(signature_end) = to_unsigned(character'pos('Z'), 8)
                then
                    audio_end_address_next <= std_ulogic_vector(u_audio_pointer + u_audio_length);
                    video_end_address_next <= std_ulogic_vector(u_audio_pointer + u_audio_length + u_video_length);

                    -- Set the pointers up to point to the 1st entry regardless of it is available or not.
                    -- This is necessary so we can check whether we are at the end of the data.
                    audio_pointer_next <= std_ulogic_vector(u_audio_pointer);
                    video_pointer_next <= std_ulogic_vector(u_audio_pointer + u_audio_length);

                    if u_audio_length /= 0 then
                        state_next <= WAIT_FOR_DATA;
                        read_audio_n_video_next <= '1';

                        memory_driver_start <= '1';
                        memory_driver_address <= audio_pointer;

                        audio_pointer_next <= std_ulogic_vector(u_audio_pointer + 1);
                    elsif u_video_length /= 0 then
                        state_next <= WAIT_FOR_DATA;
                        read_audio_n_video_next <= '0';

                        -- audio_length / video_length are only valid in PARSE_HEADER that's why we need to
                        -- calculate the address here, otherwise we would have read it from video_pointer directly.

                        memory_driver_start <= '1';
                        memory_driver_address <= std_ulogic_vector(u_audio_pointer + u_audio_length);

                        video_pointer_next <= std_ulogic_vector(u_audio_pointer + u_audio_length + 1);
                    else
                        state_next <= IDLE;
                    end if;
                else
                    state_next <= IDLE;
                    report "No media file found in memory." severity failure;
                end if;

            when WAIT_FOR_DATA =>
                if memory_driver_done = '1' then
                    state_next <= REQUEST_DATA;

                    read_audio_n_video_next <= not read_audio_n_video;

                    if read_audio_n_video = '1' then
                        audio_fifo_write_enable <= '1';

                        -- Reverse the bit order going into the Fifo because
                        -- the output is only one bit and it outputs MSB first.
                        audio_fifo_data_in <=
                            memory_driver_data(0) &
                            memory_driver_data(1) &
                            memory_driver_data(2) &
                            memory_driver_data(3) &
                            memory_driver_data(4) &
                            memory_driver_data(5) &
                            memory_driver_data(6) &
                            memory_driver_data(7)
                        ;
                    else
                        video_fifo_write_enable <= '1';

                        video_fifo_data_in <=
                            memory_driver_data(0) &
                            memory_driver_data(1) &
                            memory_driver_data(2) &
                            memory_driver_data(3) &
                            memory_driver_data(4) &
                            memory_driver_data(5) &
                            memory_driver_data(6) &
                            memory_driver_data(7)
                        ;
                    end if;
                end if;

            when REQUEST_DATA =>
                if audio_pointer = audio_end_address and video_pointer = video_end_address then
                    state_next <= DONE;

                    audio_loaded_next <= '1';
                    video_loaded_next <= '1';

                    -- We have to start playback if the audio and video data completely fit inside
                    -- the Fifos before hitting WAIT_FOR_EMPTY_SLOT.
                    if start_playback = '0' then
                        start_playback_next <= '1';

                        audio_driver_play <= '1';
                        video_driver_play <= '1';
                    end if;
                elsif read_audio_n_video = '1' then
                    if audio_fifo_full = '0' then
                        -- We are done reading audio.
                        -- Comparing two different length ulogic vector will yield false
                        -- if they are not equally long even if they are numerically the same.
                        -- Either compare as unsigned or extend to bigger vector.
                        if u_audio_pointer = unsigned(audio_end_address) then
                            read_audio_n_video_next <= '0';
                            audio_loaded_next <= '1';

                            if video_loaded = '1' then
                                start_playback_next <= '1';
                                audio_driver_play <= '1';
                                video_driver_play <= '1';
                            end if;
                        else
                            memory_driver_start <= '1';
                            memory_driver_address <= audio_pointer;

                            audio_pointer_next <= std_ulogic_vector(u_audio_pointer + 1);
                            state_next <= WAIT_FOR_DATA;
                        end if;
                    else
                        audio_loaded_next <= '1';
                        read_audio_n_video_next <= '0';
                        if video_fifo_full = '1' then
                            state_next <= WAIT_FOR_EMPTY_SLOT;
                        end if;
                    end if;
                else
                    if video_fifo_full = '0' then
                        if u_video_pointer = unsigned(video_end_address) then
                            read_audio_n_video_next <= '1';
                            video_loaded_next <= '1';

                            if audio_loaded = '1' then
                                start_playback_next <= '1';
                                audio_driver_play <= '1';
                                video_driver_play <= '1';
                            end if;
                        else
                            memory_driver_start <= '1';
                            memory_driver_address <= video_pointer;

                            video_pointer_next <= std_ulogic_vector(u_video_pointer + 1);
                            state_next <= WAIT_FOR_DATA;
                        end if;
                    else
                        video_loaded_next <= '1';
                        read_audio_n_video_next <= '1';
                        if audio_fifo_full = '1' then
                            state_next <= WAIT_FOR_EMPTY_SLOT;
                        end if;
                    end if;
                end if;

            when WAIT_FOR_EMPTY_SLOT =>
                -- If we filled both FIFOs then we can start playback
                -- incase we didn't fill both Fifos and didn't enter this stae
                -- playback starts from READ_DATA.
                if start_playback = '0' then
                    start_playback_next <= '1';

                    audio_driver_play <= '1';
                    video_driver_play <= '1';
                end if;

                if audio_fifo_full = '0' then
                    state_next <= REQUEST_DATA;
                    read_audio_n_video_next <= '1';
                elsif video_fifo_full = '0' then
                    state_next <= REQUEST_DATA;
                    read_audio_n_video_next <= '0';
                end if;

            when DONE =>
                if audio_driver_done = '1' and video_driver_done = '1' then
                    state_next <= IDLE;
                end if;
        end case;
    end process;
end architecture;
