library ieee;
use ieee.std_logic_1164.all;

entity small_led_board_tb is
end entity;

architecture tb of small_led_board_tb is

begin

end architecture;
